module avg_mag (
    input signed [17:0] decision_variable,
    input sym_clk_en, clr_acc, 
    output 
)