module GSM_filt #(
    parameter WIDTH=18,
    parameter SUM1WID=11,
    parameter SUM2WID=6,
    parameter SUM3WID=3,
    parameter SUM4WID=1
)
(

);


endmodule
