module avg_err #(parameter LFSR_WID = 22,parameter ACC_WID = 40)( 
    input signed [17:0] dec_var,
    input sym_clk_en, clr_acc, clk, reset, 
    output reg signed [17:0] ref_lvl, map_out_pwr
);

endmodule
